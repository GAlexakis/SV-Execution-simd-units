module tb;
    mul_test test ();
endmodule